* C:\Users\abyan\Documents\UT-951\ELECII\project\project2\Schematic1.sch

* Schematics Version 9.2
* Tue Jan 03 17:00:03 2017



** Analysis setup **
.tran 0ns 2m
.four 1k 5 v([$N_0001])
.OP 
.LIB "C:\Users\abyan\Documents\UT-951\ELECII\project\project2\Schematic1.lib"


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Schematic1.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
